//Files: pc.v
//Function: This block has 2 functions (1) Increase the current pc by 4 (2) Update the value of the current pc with the following pc ( I.e pc+4) or with the pc obtained from a control instruction (BEQ or JUMP). The zero flag from the ALU is used to make this decision.
//Inputs:
//clk: System clock
//arst_n: Asynchronous Reset
//enable: External signal that enables the updating of the pc when it is asserted. 
//branch_pc: Address of the branch target previously processed.
//Jump_pc: Address of the jump target previously processed.
//Zero_flag: Output of the ALU that informs if the result of the last operation is 0. This is used for processing the BEQ instructions where a subtraction between 2 operands allows to check if the condition is met.
//Branch: Signal generated by the control unit if a branch instruction is being processed.
//Jump: Signal generated by the control unit if a jump instruction is being processed.
//Outputs:
//updated_pc: Next PC used for the next clock cycle. 
//current_pc: PC that is currently processed. 


module pc#(
	parameter integer DATA_W = 16
	)(
		input  wire              clk,
		input  wire              arst_n,
		input wire              hazard,
		input  wire              enable,
		input  wire [DATA_W-1:0] branch_pc,
		input  wire [DATA_W-1:0] jump_pc,  
		input  wire              zero_flag,
		input  wire              branch,
		input  wire              jump,
		output reg  [DATA_W-1:0] updated_pc,
		output reg  [DATA_W-1:0] current_pc,
		output reg was_taken
	);

	localparam  [DATA_W-1:0] PC_INCREASE= {{(DATA_W-3){1'b0}},3'd4};

	wire [DATA_W-1:0] pc_r,next_pc,next_pc_i;
	reg               pc_src, was_taken;

	always@(*) pc_src = zero_flag & branch;
	always@(*) was_taken = zero_flag & branch;

	mux_2#(
		.DATA_W(DATA_W)
	) mux_branch( 
		.input_a (branch_pc ),
		.input_b (updated_pc),
		.select_a(pc_src    ),
		.mux_out (next_pc_i )
	);
	
	mux_2#(
		.DATA_W(DATA_W)
	) mux_jump( 
		.input_a (jump_pc   ),
		.input_b (next_pc_i ),
		.select_a(jump      ),
		.mux_out (next_pc   )
	);
	
	reg_arstn_en_hazards#(
		.DATA_W(DATA_W),
		.PRESET_VAL('b0)
	) pc_register(
		.clk   (clk       ),
		.arst_n(arst_n		),
		.hazard(hazard		),
		.din   (next_pc   ),
		.en    (enable    ),
		.dout  (current_pc)
	);

	always@(*) begin
		updated_pc = current_pc+PC_INCREASE;
	end
endmodule


